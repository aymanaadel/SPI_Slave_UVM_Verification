module spi_wrapper_sva(spi_wrapper_if.DUT s_if);
	
	// Add your Assertions here...

endmodule